-- Nandland tutorial 2
-- Joey 07Jun2020
